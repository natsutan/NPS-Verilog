module NPS_rom # (parameter DATA_WIDTH = 24 ,  ADR_WIDTH = 9)
  (
    input 			clk,
    input 			reset_x,
    input 			start,
    input 			set,
    input 			vi,
    input 			fi,
    input [ADR_WIDTH-1:0] 	datai,   
    output reg 			vo,
    output reg 			fo,
    output reg [DATA_WIDTH-1:0] datao

   );
  
  always @(posedge clk or negedge reset_x)begin
    if(reset_x == 1'b0)begin
      datao <= 0;
    end else begin
      case(datai)
	0:datao <= 24'hffffcb;
	1:datao <= 24'hfffe39;
	2:datao <= 24'hfffca8;
	3:datao <= 24'hfffb16;
	4:datao <= 24'hfff984;
	5:datao <= 24'hfff7f3;
	6:datao <= 24'hfff662;
	7:datao <= 24'hfff4d2;
	8:datao <= 24'hfff341;
	9:datao <= 24'hfff1b2;
	10:datao <= 24'hfff023;
	11:datao <= 24'hffee94;
	12:datao <= 24'hffed06;
	13:datao <= 24'hffeb79;
	14:datao <= 24'hffe9ed;
	15:datao <= 24'hffe861;
	16:datao <= 24'hffe6d7;
	17:datao <= 24'hffe54d;
	18:datao <= 24'hffe3c5;
	19:datao <= 24'hffe23d;
	20:datao <= 24'hffe0b7;
	21:datao <= 24'hffdf32;
	22:datao <= 24'hffddae;
	23:datao <= 24'hffdc2b;
	24:datao <= 24'hffdaaa;
	25:datao <= 24'hffd92a;
	26:datao <= 24'hffd7ac;
	27:datao <= 24'hffd630;
	28:datao <= 24'hffd4b5;
	29:datao <= 24'hffd33b;
	30:datao <= 24'hffd1c3;
	31:datao <= 24'hffd04e;
	32:datao <= 24'hffceda;
	33:datao <= 24'hffcd67;
	34:datao <= 24'hffcbf7;
	35:datao <= 24'hffca89;
	36:datao <= 24'hffc91d;
	37:datao <= 24'hffc7b3;
	38:datao <= 24'hffc64b;
	39:datao <= 24'hffc4e5;
	40:datao <= 24'hffc382;
	41:datao <= 24'hffc221;
	42:datao <= 24'hffc0c2;
	43:datao <= 24'hffbf66;
	44:datao <= 24'hffbe0c;
	45:datao <= 24'hffbcb5;
	46:datao <= 24'hffbb61;
	47:datao <= 24'hffba0f;
	48:datao <= 24'hffb8bf;
	49:datao <= 24'hffb773;
	50:datao <= 24'hffb629;
	51:datao <= 24'hffb4e2;
	52:datao <= 24'hffb39e;
	53:datao <= 24'hffb25d;
	54:datao <= 24'hffb11f;
	55:datao <= 24'hffafe4;
	56:datao <= 24'hffaeac;
	57:datao <= 24'hffad77;
	58:datao <= 24'hffac46;
	59:datao <= 24'hffab17;
	60:datao <= 24'hffa9ec;
	61:datao <= 24'hffa8c4;
	62:datao <= 24'hffa7a0;
	63:datao <= 24'hffa67f;
	64:datao <= 24'hffa561;
	65:datao <= 24'hffa447;
	66:datao <= 24'hffa331;
	67:datao <= 24'hffa21e;
	68:datao <= 24'hffa10e;
	69:datao <= 24'hffa003;
	70:datao <= 24'hff9efb;
	71:datao <= 24'hff9df6;
	72:datao <= 24'hff9cf6;
	73:datao <= 24'hff9bf9;
	74:datao <= 24'hff9b00;
	75:datao <= 24'hff9a0b;
	76:datao <= 24'hff991a;
	77:datao <= 24'hff982d;
	78:datao <= 24'hff9744;
	79:datao <= 24'hff965f;
	80:datao <= 24'hff957e;
	81:datao <= 24'hff94a1;
	82:datao <= 24'hff93c8;
	83:datao <= 24'hff92f4;
	84:datao <= 24'hff9223;
	85:datao <= 24'hff9157;
	86:datao <= 24'hff908f;
	87:datao <= 24'hff8fcc;
	88:datao <= 24'hff8f0d;
	89:datao <= 24'hff8e52;
	90:datao <= 24'hff8d9b;
	91:datao <= 24'hff8ce9;
	92:datao <= 24'hff8c3b;
	93:datao <= 24'hff8b92;
	94:datao <= 24'hff8aed;
	95:datao <= 24'hff8a4d;
	96:datao <= 24'hff89b1;
	97:datao <= 24'hff891a;
	98:datao <= 24'hff8888;
	99:datao <= 24'hff87fa;
	100:datao <= 24'hff8770;
	101:datao <= 24'hff86ec;
	102:datao <= 24'hff866c;
	103:datao <= 24'hff85f0;
	104:datao <= 24'hff8579;
	105:datao <= 24'hff8508;
	106:datao <= 24'hff849a;
	107:datao <= 24'hff8432;
	108:datao <= 24'hff83ce;
	109:datao <= 24'hff836f;
	110:datao <= 24'hff8315;
	111:datao <= 24'hff82c0;
	112:datao <= 24'hff826f;
	113:datao <= 24'hff8224;
	114:datao <= 24'hff81dd;
	115:datao <= 24'hff819b;
	116:datao <= 24'hff815e;
	117:datao <= 24'hff8126;
	118:datao <= 24'hff80f2;
	119:datao <= 24'hff80c4;
	120:datao <= 24'hff809b;
	121:datao <= 24'hff8076;
	122:datao <= 24'hff8056;
	123:datao <= 24'hff803c;
	124:datao <= 24'hff8026;
	125:datao <= 24'hff8015;
	126:datao <= 24'hff8009;
	127:datao <= 24'hff8002;
	128:datao <= 24'hff8000;
	129:datao <= 24'hff8002;
	130:datao <= 24'hff800a;
	131:datao <= 24'hff8017;
	132:datao <= 24'hff8028;
	133:datao <= 24'hff803f;
	134:datao <= 24'hff805a;
	135:datao <= 24'hff807a;
	136:datao <= 24'hff80a0;
	137:datao <= 24'hff80ca;
	138:datao <= 24'hff80f9;
	139:datao <= 24'hff812d;
	140:datao <= 24'hff8166;
	141:datao <= 24'hff81a3;
	142:datao <= 24'hff81e6;
	143:datao <= 24'hff822d;
	144:datao <= 24'hff827a;
	145:datao <= 24'hff82cb;
	146:datao <= 24'hff8321;
	147:datao <= 24'hff837b;
	148:datao <= 24'hff83db;
	149:datao <= 24'hff843f;
	150:datao <= 24'hff84a8;
	151:datao <= 24'hff8516;
	152:datao <= 24'hff8589;
	153:datao <= 24'hff8600;
	154:datao <= 24'hff867c;
	155:datao <= 24'hff86fd;
	156:datao <= 24'hff8782;
	157:datao <= 24'hff880c;
	158:datao <= 24'hff889a;
	159:datao <= 24'hff892e;
	160:datao <= 24'hff89c5;
	161:datao <= 24'hff8a62;
	162:datao <= 24'hff8b02;
	163:datao <= 24'hff8ba8;
	164:datao <= 24'hff8c52;
	165:datao <= 24'hff8d00;
	166:datao <= 24'hff8db3;
	167:datao <= 24'hff8e6a;
	168:datao <= 24'hff8f25;
	169:datao <= 24'hff8fe5;
	170:datao <= 24'hff90a9;
	171:datao <= 24'hff9172;
	172:datao <= 24'hff923e;
	173:datao <= 24'hff930f;
	174:datao <= 24'hff93e4;
	175:datao <= 24'hff94be;
	176:datao <= 24'hff959b;
	177:datao <= 24'hff967c;
	178:datao <= 24'hff9762;
	179:datao <= 24'hff984c;
	180:datao <= 24'hff9939;
	181:datao <= 24'hff9a2b;
	182:datao <= 24'hff9b20;
	183:datao <= 24'hff9c1a;
	184:datao <= 24'hff9d17;
	185:datao <= 24'hff9e18;
	186:datao <= 24'hff9f1d;
	187:datao <= 24'hffa025;
	188:datao <= 24'hffa131;
	189:datao <= 24'hffa241;
	190:datao <= 24'hffa355;
	191:datao <= 24'hffa46c;
	192:datao <= 24'hffa586;
	193:datao <= 24'hffa6a4;
	194:datao <= 24'hffa7c6;
	195:datao <= 24'hffa8eb;
	196:datao <= 24'hffaa13;
	197:datao <= 24'hffab3e;
	198:datao <= 24'hffac6d;
	199:datao <= 24'hffad9f;
	200:datao <= 24'hffaed5;
	201:datao <= 24'hffb00d;
	202:datao <= 24'hffb148;
	203:datao <= 24'hffb287;
	204:datao <= 24'hffb3c8;
	205:datao <= 24'hffb50d;
	206:datao <= 24'hffb654;
	207:datao <= 24'hffb79e;
	208:datao <= 24'hffb8eb;
	209:datao <= 24'hffba3a;
	210:datao <= 24'hffbb8d;
	211:datao <= 24'hffbce2;
	212:datao <= 24'hffbe39;
	213:datao <= 24'hffbf93;
	214:datao <= 24'hffc0f0;
	215:datao <= 24'hffc24f;
	216:datao <= 24'hffc3b0;
	217:datao <= 24'hffc514;
	218:datao <= 24'hffc67a;
	219:datao <= 24'hffc7e2;
	220:datao <= 24'hffc94c;
	221:datao <= 24'hffcab8;
	222:datao <= 24'hffcc27;
	223:datao <= 24'hffcd97;
	224:datao <= 24'hffcf0a;
	225:datao <= 24'hffd07e;
	226:datao <= 24'hffd1f4;
	227:datao <= 24'hffd36c;
	228:datao <= 24'hffd4e6;
	229:datao <= 24'hffd661;
	230:datao <= 24'hffd7de;
	231:datao <= 24'hffd95c;
	232:datao <= 24'hffdadc;
	233:datao <= 24'hffdc5d;
	234:datao <= 24'hffdde0;
	235:datao <= 24'hffdf64;
	236:datao <= 24'hffe0e9;
	237:datao <= 24'hffe270;
	238:datao <= 24'hffe3f8;
	239:datao <= 24'hffe580;
	240:datao <= 24'hffe70a;
	241:datao <= 24'hffe895;
	242:datao <= 24'hffea20;
	243:datao <= 24'hffebad;
	244:datao <= 24'hffed3a;
	245:datao <= 24'hffeec8;
	246:datao <= 24'hfff056;
	247:datao <= 24'hfff1e6;
	248:datao <= 24'hfff375;
	249:datao <= 24'hfff506;
	250:datao <= 24'hfff696;
	251:datao <= 24'hfff827;
	252:datao <= 24'hfff9b8;
	253:datao <= 24'hfffb4a;
	254:datao <= 24'hfffcdc;
	255:datao <= 24'hfffe6e;
	256:datao <= 24'h0;
	257:datao <= 24'h191;
	258:datao <= 24'h323;
	259:datao <= 24'h4b5;
	260:datao <= 24'h647;
	261:datao <= 24'h7d8;
	262:datao <= 24'h969;
	263:datao <= 24'haf9;
	264:datao <= 24'hc8a;
	265:datao <= 24'he19;
	266:datao <= 24'hfa9;
	267:datao <= 24'h1137;
	268:datao <= 24'h12c5;
	269:datao <= 24'h1452;
	270:datao <= 24'h15df;
	271:datao <= 24'h176a;
	272:datao <= 24'h18f5;
	273:datao <= 24'h1a7f;
	274:datao <= 24'h1c07;
	275:datao <= 24'h1d8f;
	276:datao <= 24'h1f16;
	277:datao <= 24'h209b;
	278:datao <= 24'h221f;
	279:datao <= 24'h23a2;
	280:datao <= 24'h2523;
	281:datao <= 24'h26a3;
	282:datao <= 24'h2821;
	283:datao <= 24'h299e;
	284:datao <= 24'h2b19;
	285:datao <= 24'h2c93;
	286:datao <= 24'h2e0b;
	287:datao <= 24'h2f81;
	288:datao <= 24'h30f5;
	289:datao <= 24'h3268;
	290:datao <= 24'h33d8;
	291:datao <= 24'h3547;
	292:datao <= 24'h36b3;
	293:datao <= 24'h381d;
	294:datao <= 24'h3985;
	295:datao <= 24'h3aeb;
	296:datao <= 24'h3c4f;
	297:datao <= 24'h3db0;
	298:datao <= 24'h3f0f;
	299:datao <= 24'h406c;
	300:datao <= 24'h41c6;
	301:datao <= 24'h431d;
	302:datao <= 24'h4472;
	303:datao <= 24'h45c5;
	304:datao <= 24'h4714;
	305:datao <= 24'h4861;
	306:datao <= 24'h49ab;
	307:datao <= 24'h4af2;
	308:datao <= 24'h4c37;
	309:datao <= 24'h4d78;
	310:datao <= 24'h4eb7;
	311:datao <= 24'h4ff2;
	312:datao <= 24'h512a;
	313:datao <= 24'h5260;
	314:datao <= 24'h5392;
	315:datao <= 24'h54c1;
	316:datao <= 24'h55ec;
	317:datao <= 24'h5714;
	318:datao <= 24'h5839;
	319:datao <= 24'h595b;
	320:datao <= 24'h5a79;
	321:datao <= 24'h5b93;
	322:datao <= 24'h5caa;
	323:datao <= 24'h5dbe;
	324:datao <= 24'h5ece;
	325:datao <= 24'h5fda;
	326:datao <= 24'h60e2;
	327:datao <= 24'h61e7;
	328:datao <= 24'h62e8;
	329:datao <= 24'h63e5;
	330:datao <= 24'h64df;
	331:datao <= 24'h65d4;
	332:datao <= 24'h66c6;
	333:datao <= 24'h67b3;
	334:datao <= 24'h689d;
	335:datao <= 24'h6983;
	336:datao <= 24'h6a64;
	337:datao <= 24'h6b41;
	338:datao <= 24'h6c1b;
	339:datao <= 24'h6cf0;
	340:datao <= 24'h6dc1;
	341:datao <= 24'h6e8d;
	342:datao <= 24'h6f56;
	343:datao <= 24'h701a;
	344:datao <= 24'h70da;
	345:datao <= 24'h7195;
	346:datao <= 24'h724c;
	347:datao <= 24'h72ff;
	348:datao <= 24'h73ad;
	349:datao <= 24'h7457;
	350:datao <= 24'h74fd;
	351:datao <= 24'h759d;
	352:datao <= 24'h763a;
	353:datao <= 24'h76d1;
	354:datao <= 24'h7765;
	355:datao <= 24'h77f3;
	356:datao <= 24'h787d;
	357:datao <= 24'h7902;
	358:datao <= 24'h7983;
	359:datao <= 24'h79ff;
	360:datao <= 24'h7a76;
	361:datao <= 24'h7ae9;
	362:datao <= 24'h7b57;
	363:datao <= 24'h7bc0;
	364:datao <= 24'h7c24;
	365:datao <= 24'h7c84;
	366:datao <= 24'h7cde;
	367:datao <= 24'h7d34;
	368:datao <= 24'h7d85;
	369:datao <= 24'h7dd2;
	370:datao <= 24'h7e19;
	371:datao <= 24'h7e5c;
	372:datao <= 24'h7e99;
	373:datao <= 24'h7ed2;
	374:datao <= 24'h7f06;
	375:datao <= 24'h7f35;
	376:datao <= 24'h7f5f;
	377:datao <= 24'h7f85;
	378:datao <= 24'h7fa5;
	379:datao <= 24'h7fc0;
	380:datao <= 24'h7fd7;
	381:datao <= 24'h7fe8;
	382:datao <= 24'h7ff5;
	383:datao <= 24'h7ffd;
	384:datao <= 24'h7fff;
	385:datao <= 24'h7ffd;
	386:datao <= 24'h7ff6;
	387:datao <= 24'h7fea;
	388:datao <= 24'h7fd9;
	389:datao <= 24'h7fc3;
	390:datao <= 24'h7fa9;
	391:datao <= 24'h7f89;
	392:datao <= 24'h7f64;
	393:datao <= 24'h7f3b;
	394:datao <= 24'h7f0d;
	395:datao <= 24'h7ed9;
	396:datao <= 24'h7ea1;
	397:datao <= 24'h7e64;
	398:datao <= 24'h7e22;
	399:datao <= 24'h7ddb;
	400:datao <= 24'h7d90;
	401:datao <= 24'h7d3f;
	402:datao <= 24'h7cea;
	403:datao <= 24'h7c90;
	404:datao <= 24'h7c31;
	405:datao <= 24'h7bcd;
	406:datao <= 24'h7b65;
	407:datao <= 24'h7af7;
	408:datao <= 24'h7a86;
	409:datao <= 24'h7a0f;
	410:datao <= 24'h7993;
	411:datao <= 24'h7913;
	412:datao <= 24'h788f;
	413:datao <= 24'h7805;
	414:datao <= 24'h7777;
	415:datao <= 24'h76e5;
	416:datao <= 24'h764e;
	417:datao <= 24'h75b2;
	418:datao <= 24'h7512;
	419:datao <= 24'h746d;
	420:datao <= 24'h73c4;
	421:datao <= 24'h7316;
	422:datao <= 24'h7264;
	423:datao <= 24'h71ad;
	424:datao <= 24'h70f2;
	425:datao <= 24'h7033;
	426:datao <= 24'h6f70;
	427:datao <= 24'h6ea8;
	428:datao <= 24'h6ddc;
	429:datao <= 24'h6d0b;
	430:datao <= 24'h6c37;
	431:datao <= 24'h6b5e;
	432:datao <= 24'h6a81;
	433:datao <= 24'h69a0;
	434:datao <= 24'h68bb;
	435:datao <= 24'h67d2;
	436:datao <= 24'h66e5;
	437:datao <= 24'h65f4;
	438:datao <= 24'h64ff;
	439:datao <= 24'h6406;
	440:datao <= 24'h6309;
	441:datao <= 24'h6209;
	442:datao <= 24'h6104;
	443:datao <= 24'h5ffc;
	444:datao <= 24'h5ef1;
	445:datao <= 24'h5de1;
	446:datao <= 24'h5cce;
	447:datao <= 24'h5bb8;
	448:datao <= 24'h5a9e;
	449:datao <= 24'h5980;
	450:datao <= 24'h585f;
	451:datao <= 24'h573b;
	452:datao <= 24'h5613;
	453:datao <= 24'h54e8;
	454:datao <= 24'h53b9;
	455:datao <= 24'h5288;
	456:datao <= 24'h5153;
	457:datao <= 24'h501b;
	458:datao <= 24'h4ee0;
	459:datao <= 24'h4da2;
	460:datao <= 24'h4c61;
	461:datao <= 24'h4b1d;
	462:datao <= 24'h49d6;
	463:datao <= 24'h488c;
	464:datao <= 24'h4740;
	465:datao <= 24'h45f0;
	466:datao <= 24'h449e;
	467:datao <= 24'h434a;
	468:datao <= 24'h41f3;
	469:datao <= 24'h4099;
	470:datao <= 24'h3f3d;
	471:datao <= 24'h3dde;
	472:datao <= 24'h3c7d;
	473:datao <= 24'h3b1a;
	474:datao <= 24'h39b4;
	475:datao <= 24'h384c;
	476:datao <= 24'h36e2;
	477:datao <= 24'h3576;
	478:datao <= 24'h3408;
	479:datao <= 24'h3298;
	480:datao <= 24'h3125;
	481:datao <= 24'h2fb1;
	482:datao <= 24'h2e3c;
	483:datao <= 24'h2cc4;
	484:datao <= 24'h2b4a;
	485:datao <= 24'h29cf;
	486:datao <= 24'h2853;
	487:datao <= 24'h26d5;
	488:datao <= 24'h2555;
	489:datao <= 24'h23d4;
	490:datao <= 24'h2251;
	491:datao <= 24'h20cd;
	492:datao <= 24'h1f48;
	493:datao <= 24'h1dc2;
	494:datao <= 24'h1c3a;
	495:datao <= 24'h1ab2;
	496:datao <= 24'h1928;
	497:datao <= 24'h179e;
	498:datao <= 24'h1612;
	499:datao <= 24'h1486;
	500:datao <= 24'h12f9;
	501:datao <= 24'h116b;
	502:datao <= 24'hfdc;
	503:datao <= 24'he4d;
	504:datao <= 24'hcbe;
	505:datao <= 24'hb2d;
	506:datao <= 24'h99d;
	507:datao <= 24'h80c;
	508:datao <= 24'h67b;
	509:datao <= 24'h4e9;
	510:datao <= 24'h357;
	511:datao <= 24'h1c6;
      endcase
    end
  end // always @ (posedge clk or negedge reset_x)
  

  always @ (posedge clk or negedge reset_x) begin
    if(reset_x == 1'b0)begin
      vo <= 0;
      fo <= 0;
    end else begin
      vo <= vi;
      fo <= fi;
    end
  end
  
  

  
endmodule
